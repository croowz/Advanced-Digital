`timescale 1ns/1ps

module toy_tbw_tb_0;

	reg CLK = 1'b0;
	reg [7:0] D_IN = 8'b00000000;
	reg RESET = 1'b1; 

	wire [7:0] ADDR; 	
	wire [7:0] D_OUT; 
	wire MEM_EN;
	wire RORW; 
	wire S0;
	wire S1;
	wire S2;
	wire S3; 
	wire S4; 
	wire S5;

	initial // Clock process for CLK 
		begin 
			forever 
				begin
					CLK = 1'b0;
					#50; 
					CLK = 1'b1; 
					#50;
				end 
		end
		
	toy_sch UUT ( 
	.CLK(CLK), 
	.D_IN(D_IN),
	.RESET(RESET),
	.ADDR(ADDR), 
	.D_OUT(D_OUT), 
	.MEM_EN(MEM_EN), 
	.RORW(RORW), 
	.S0(S0),
	.S1(S1), 
	.S2(S2), 
	.S3(S3), 
	.S4(S4), 
	.S5(S5));
	
	initial 
		begin
			// ------------- Current Time: 135ns 
			#135;
			RESET = 1'b0;
			// -------------------------------------
			
			// ------------- Current Time: 235ns 
			#100;
			D_IN = 8'b00000001;
			// -------------------------------------
			
			// ------------- Current Time: 335ns 
			#100;
			D_IN = 8'b00000000;
			// -------------------------------------
			
			// ------------- Current Time: 435ns 
			#100;
			D_IN = 8'b10101010;
			// -------------------------------------
			
			// ------------- Current Time: 535ns
			#100;
			D_IN = 8'b00000000;
			// -------------------------------------
			
			// ------------- Current Time: 735ns 
			#200;
			D_IN = 8'b00000100;
			// -------------------------------------
			
			// ------------- Current Time: 835ns 
			#100;
			D_IN = 8'b00000000;
			// -------------------------------------
			
			// ------------- Current Time: 1035ns 
			#200;
			D_IN = 8'b00000001;
			// -------------------------------------
			
			// ------------- Current Time: 1135ns 
			#100;
			D_IN = 8'b00000000;
			// -------------------------------------
			
			// ------------- Current Time: 1235ns 
			#100;
			D_IN = 8'b11111110;
			// -------------------------------------
			
			// ------------- Current Time: 1335ns 
			#100;
			D_IN = 8'b00000000;
			// -------------------------------------
			
			// ------------- Current Time: 1535ns 
			#200;
			D_IN = 8'b00000010;
			// -------------------------------------
			
			// ------------- Current Time: 1635ns 
			#100;
			D_IN = 8'b00000000;
			// -------------------------------------
			
			// ------------- Current Time: 1735ns 
			#100;
			D_IN = 8'b00000011;/////*********
			// -------------------------------------
			
			// ------------- Current Time: 1835ns 
			#100;
			D_IN = 8'b00000000;
			// -------------------------------------
			
			// ------------- Current Time: 2035ns 
			#200;
			D_IN = 8'b00010000;
			// -------------------------------------
			
			// ------------- Current Time: 2135ns 
			#100;
			D_IN = 8'b00000000;
			// -------------------------------------
			
			// ------------- Current Time: 2235ns 
			#100;
			D_IN = 8'b11111111;
			// -------------------------------------
			
			// ------------- Current Time: 2335ns 
			#100;
			D_IN = 8'b00000000;
			// -------------------------------------
			
			// ------------- Current Time: 2535ns 
			#200;
			D_IN = 8'b00000100;
			// -------------------------------------
			
			// ------------- Current Time: 2635ns 
			#100;
			D_IN = 8'b00000000;
			// -------------------------------------
			
			// ------------- Current Time: 2835ns 
			#200;
			D_IN = 8'b00001000;
			// -------------------------------------
			
			// ------------- Current Time: 2935ns 
			#100;
			D_IN = 8'b00000000;
			// -------------------------------------
			
			// ------------- Current Time: 3035ns 
			#100;
			D_IN = 8'b11001100;
			// -------------------------------------
			
			// ------------- Current Time: 3135ns 
			#100;
			D_IN = 8'b00000000;
			// -------------------------------------
			
			// ------------- Current Time: 3335ns 
			#200;
			D_IN = 8'b00000001;
			// -------------------------------------
			
			// ------------- Current Time: 3435ns 
			#100;
			D_IN = 8'b00000000;
			// -------------------------------------
			
			// ------------- Current Time: 3535ns 
			#100;
			D_IN = 8'b00001111;
			// -------------------------------------
			
			// ------------- Current Time: 3635ns 
			#100;
			D_IN = 8'b00000000;
			// -------------------------------------
			
			// ------------- Current Time: 3835ns 
			#200;
			D_IN = 8'b00001000;
			// -------------------------------------
			
			// ------------- Current Time: 3935ns 
			#100;
			D_IN = 8'b00000000;
			// -------------------------------------
			
			// ------------- Current Time: 4035ns 
			#100;
			D_IN = 8'b11111110;
			// -------------------------------------
			
			// ------------- Current Time: 4135ns 
			#100;
			D_IN = 8'b00000000;
			// -------------------------------------
		end 
endmodule
