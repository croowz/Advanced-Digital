`timescale 1ns/1ps

module mux8_tbw_tb_0;
	reg [7:0] IN0 = 8'b00000000;
	reg [7:0] IN1 = 8'b00000000;
	reg SEL = 1'b0;

	wire [7:0] MUX_OUT;

	mux8sch UUT (
		.IN0(IN0),
		.IN1(IN1),
		.SEL(SEL),
		.MUX_OUT(MUX_OUT));

	initial 
		begin
			// ------------- Current Time: 100ns
			#100;
			IN1 = 8'b01011111;
			// -------------------------------------
			
			// ------------- Current Time: 200ns
			#100;
			SEL = 1'b1;
			IN0 = 8'b01011111;
			IN1 = 8'b11001000;
			// -------------------------------------
			
			// ------------- Current Time: 300ns
			#100;
			IN1 = 8'b10010001;
			// -------------------------------------
			
			// ------------- Current Time: 400ns
			#100;
			IN0 = 8'b11001000;
			IN1 = 8'b00011101;
			// -------------------------------------
			
			// ------------- Current Time: 500ns
			#100;
			SEL = 1'b0;
			IN1 = 8'b11101010;
			// -------------------------------------
			
			// ------------- Current Time: 600ns
			#100;
			IN0 = 8'b10010001;
			IN1 = 8'b01110011;
			// -------------------------------------
			
			// ------------- Current Time: 700ns
			#100;
			SEL = 1'b1;
			IN1 = 8'b01110100;
			// -------------------------------------
			
			// ------------- Current Time: 800ns
			#100;
			IN0 = 8'b00011101;
			IN1 = 8'b10101000;
			// -------------------------------------
			
			// ------------- Current Time: 1000ns
			#200;
			IN0 = 8'b11101010;
			//--------------------------------------
		end
endmodule
