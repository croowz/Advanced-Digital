/*
 * Design: CSEE4270 - Skeleton Module for Binary to BCD Converter
 * Author: 
 * 
 *
 * 
 *
 */

`timescale 1ns / 1ns
module Binary2BCD(Cnt, Tens, Ones);

   input [3:0] Cnt;
   output [3:0] Tens, Ones;

endmodule
